module Connection_ports_by_name ( input a, input b, output out );
    mod_a test(.out(out),.in1(a),.in2(b));
endmodule
