module modules ( input a, input b, output out );
    mod_a test(.out(out),.in1(a),.in2(b));
endmodule